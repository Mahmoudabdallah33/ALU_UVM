package pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "ALU_seq_item.sv"
`include "ALU_sqr.sv"
`include "agt_config.sv"
`include "env_config.sv"
`include "ALU_seq.sv"
`include "ALU_vseq.sv"
`include "ALU_drv.sv"
`include "ALU_mon.sv"
`include "ALU_agt.sv"
`include "ALU_evaluator.sv"
`include "ALU_predictor.sv"
`include "ALU_scb.sv"
`include "ALU_cov.sv"
`include "ALU_env.sv"
`include "ALU_test.sv"




endpackage

